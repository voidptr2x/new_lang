module v_backend

pub fn bprint(str string, nline string)
{
	
}