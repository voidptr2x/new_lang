module parser

pub fn (mut b B_Lang) parse_struct(struct_code []string) string {
	return ""
}